module ysyx_22041412_if(
    input clk,
    input rst,
//performance counter
    output reg [63:0]       pred_miss_count,
    output reg [63:0]       pred_hit_count,

    output reg[63:0]pc,
    output reg[31:0]imm_data,

    input jarl_rady,
    input valid_i,  //ID OK
    output reg ready_o,  

    //跳转处理部分
    //跳转处理部分
    //input   jump_hit,          //1 分支结果为跳转   0不跳    为分支预测预留的引脚
    //跳转处理部分       
    //input   jump_hit,          //1 分支结果为跳转   0不跳    为分支预测预留的引脚
    input [31:0]jal_pc,
    input       jal_ok  ,
    input       jal_b_hit,        //1 分支结果为跳转   0不跳    为分支预测使用的引脚
    input [63:0]mem_dnpc,        //其他跳转的结果

    output reg  fence_i,
    input       fence_ready,
    //ifu   <---> cache 
    input       ready_i,        // 读有效等待接收

       
    input      [31:0]r_data_i,  // 读数据
    output reg [31:0]r_addr_o,  // 读地址

    output reg if_read_vaild   //IFU读cache
 );
`define IF_IDLE         3'b000  
`define IF_WORK         3'b001 
`define IF_WAIT         3'b010 //其他跳转处理
`define IF_BRANCH       3'b100 //条件分支的处理
`define IF_FENCE        3'b111 //FENCE I

reg  [2:0] state;            //状态机 
reg  [31:0]dnpc;
//-------------快速解码部分 BEGIN----------------------
wire jump ;
wire jump_b;
wire jal ;
wire jarl;
wire ecall ;
assign fence_i  = (imm_data[6:0]==`ysyx_22041412_FENCE) ? imm_data[12] : 1'b0;
assign jal  = ( imm_data[6:0]==`ysyx_22041412_jal) ?1'b1:1'b0;  //直接跳转命令  可以直接出结果 由 译码部分计算
assign jarl = ( imm_data[6:0]==`ysyx_22041412_jalr)?1'b1:1'b0;  //直接跳转  但是需要等读取寄存器
assign ecall= (imm_data[6:0]==`ysyx_22041412_Environment & (imm_data[31:20]==12'b00000000000 || imm_data[31:20]==12'b001100000010))? 1'b1 : 1'b0;
              //ECALL MRET
assign jump_b =(imm_data[6:0]==`ysyx_22041412_B_type) ? 1'b1 : 1'b0 ;           //这段可以用分支预测
assign jump= (jump_b  | jarl | ecall ) ? 1'b1 : 1'b0;
  //针对循环的预测
    wire [31:0]B_pc  ;
    wire jump_pred   ;
    reg jump_pred_ld ;  //暂存的本次预测结果  1为直接跳  0为不跳
    assign B_pc		=	jump_b ? ( {{20{imm_data[31]}},imm_data[7],imm_data[30:25],imm_data[11:8],1'b0} + pc[31:0] ) : 32'b0;  //B类指令的目标地址
    /* 
      一条for翻译成汇编是
      xxx：
      ....
      bne loopnnum , xxx:
      如果xxx地址比当前pc小就可以认为跳，只有最后一次循环退出才会预测错一次
     */
    assign jump_pred = jump_b ? (B_pc < pc[31:0]) ?1'b1 :1'b0:1'b0;
//-------------快速解码部分 END ----------------------

    reg branch_op;
    reg branch_ok;
    reg [31:0]jump_pc;
    wire pred_hit =  (jump_pred_ld & jal_b_hit) | (~jump_pred_ld & ~jal_b_hit);
    wire pred_miss=  ~pred_hit;

    reg [31:0]pred_pc;
    reg [31:0]pred_imm;
    reg       pred_redy;

  // always @(posedge clk) begin
  //    $display("IF clk 1 oneline=%d state=%b jar %b",one_line,state,jar);
  // end  


  always@(posedge clk)begin //IFU状态机
    if(rst )begin
      state <= `IF_WORK;
    end else begin
      case (state)
        `IF_IDLE: begin
            state<= valid_i ? `IF_WORK : `IF_IDLE;
        end
        `IF_WORK:begin
            state <=(valid_i & jump ) ? `IF_WAIT 
                            : fence_i ? `IF_FENCE  : `IF_WORK;
        end
        `IF_BRANCH:begin
            state <= jarl_rady ? `IF_WORK : `IF_BRANCH;
        end
        `IF_WAIT:begin
            state <= jarl_rady ? `IF_WORK : `IF_WAIT;
        end
        `IF_FENCE:begin
            state <= fence_ready ? `IF_WORK :`IF_FENCE;
        end
        default: ;
      endcase
    end
  end

    always@(*)begin //负责转发cache的数据
        case (state)
            `IF_WORK: begin
                if (ready_i & ~last_stall)begin
                    imm_data = r_data_i;
                    pc[31:0] = r_addr_o;
                    ready_o  = 1'b1;
                end else if(last_stall)begin
                    imm_data = last_imm;
                    pc[31:0] = last_pc;
                    ready_o  = 1'b1;   
                end
                else begin
                    imm_data = 32'b0;
                    pc[31:0] = 32'b0;
                    ready_o  = 1'b0;
                end
            end
            `IF_BRANCH: begin
                if (pred_hit)begin
                    imm_data = r_data_i;
                    pc[31:0] = r_addr_o;
                    ready_o  = 1'b1;
                end else begin
                    imm_data = 32'b0;
                    pc[31:0] = 32'b0;
                    ready_o  = 1'b0;
                end
            end
            `IF_FENCE: begin
                ready_o = valid_i;
            end
            default : begin
                    imm_data = 32'b0;
                    pc[31:0] = 32'b0;
                    ready_o  = 1'b0;
            end
        endcase
    end


 reg [31:0]last_imm;
 reg [31:0]last_pc;
 reg last_stall;
 reg wait_jal;
 always @(posedge clk) begin   //IFU  DNPC控制  -->> ICACHE
  if(rst)begin
    if_read_vaild  <= 1'b1;
    dnpc           <= 32'h80000004;
    r_addr_o       <= 32'h80000000;
  end  else begin   
    case (state)
        `IF_IDLE: begin
            if_read_vaild  <= 1'b0;
            dnpc           <= dnpc;
        end
        `IF_WORK:begin
          if(~valid_i & ready_i)begin //如果发出请求后ID暂停，需要先缓存下来数据
            last_imm       <= r_data_i;
            last_pc        <= r_addr_o;
            last_stall     <= 1'b1;
            if_read_vaild  <= 1'b0;
          end 
          if(valid_i & ready_i & ~wait_jal)begin //每次取回指令后发出一条新的指令请求，地址递增+4
            if_read_vaild  <= (~jump & ~jal);
            wait_jal       <= jal;
            r_addr_o       <=dnpc;
            dnpc           <=dnpc+4;
            last_stall     <=1'b0;
            //$display("IFU Read one line : addr:%8h :%8h",dnpc,imm_data_4mux1);           
          end else if(last_stall & valid_i)begin
            if_read_vaild  <= (~jump & ~jal);
            wait_jal       <= jal;
            r_addr_o       <=dnpc;
            dnpc           <=dnpc+4;
            last_stall     <=1'b0;
          end
          else if (wait_jal & jal_ok)begin
            wait_jal       <= 1'b0;
            if_read_vaild  <= 1'b1;
            r_addr_o       <= jal_pc;
            dnpc           <= jal_pc+4;
            last_stall     <=1'b0;
          end
        //   else if(jump_b)begin
        //     if_read_vaild <= 1'b1;
        //     dnpc          <= jump_pred ? B_pc : dnpc+4 ;
        //   end

        end
        `IF_WAIT:begin       //等待分支指令给出新地址
          last_stall     <=1'b0;
          if(jarl_rady) begin
            if_read_vaild  <= 1'b1;
            r_addr_o       <= mem_dnpc[31:0];
            dnpc           <= mem_dnpc[31:0]+4;
            //$display("IFU JUMP JARL/B PC %8h",mem_dnpc[31:0]);
          end
        end
        `IF_BRANCH:begin    //条件分支的处理
            last_stall     <=1'b0;
            if(jarl_rady) begin// 结果出来了
                if(pred_hit) begin
                    pred_hit_count <= pred_hit_count+1 ;
                    //命中 直接让流水线动起来

                end
                else  begin
                    pred_miss_count <= pred_miss_count+1;
                    //MISS 需清空预取数据重新取

                end
                jump_pred_ld<= 1'b0;
            end else begin
                jump_pred_ld<= jump_pred_ld;
            end
        end
        `IF_FENCE:begin    //等待cache处理完fence
   
        end
        default: ;  
    endcase

  end

 end
endmodule
