module ysyx_22041412_i_cache(
    parameter cache_l = 'd8;
    parameter cache_line_num = 'd8;
)(

);

endmodule